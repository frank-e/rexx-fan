3��Ћ��؎���� |��� ���D�t� �VW� �� p^_����?U��k�u]����?����x�uNf�wf�D�B����r=���U��k�u2����
magic AWOL 
no boot partition 
read error ���
�t	� ����������                                                                                                                                                                                                                                                                     a5�  �                                                          U��; REXXFAT     �          � )w2�NO NAME    FAT12   �K boot code placeholder for  V�
�t	� ����^�WP��� ���P$<
i/�X��X_��  �|�|���^�����|���<�����- ���֋L�������|�����������                                                                                                                                                                                                                                                                                                       U����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             conectix      ��������� REXX  Wi2k      "       " ���   ��槹A[꺖F��PlJ�K                                                                                                                                                                                                                                                                                                                                                                                                                                            